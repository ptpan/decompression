module pip_1();








endmodule