module pip_2();






endmodule